//------------------------------------------------------------------------------
// clock_if interface
//
// This interface provides a clock output signal.
// 
//------------------------------------------------------------------------------
interface pc_if ();
    // pc output signal.
    logic[31:0] pc;
endinterface : pc_if

