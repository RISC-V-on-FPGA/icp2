//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// import uvm_pkg::*;
// `include "uvm_macros.svh"
// `include "pc_seq_item.svh"  // Include the item file

class pc_seq extends uvm_sequence #(pc_seq_item);
    `uvm_object_utils(pc_seq)

    rand bit [31:0] pc;
    int unsigned MAX_VALUE_32 = 4294967295;

    // the program count can oly be an even number
    constraint pc_c {
        pc % 2 == 0;
    }

    constraint pc_weight_c {
        pc dist { 0              :/ 2, 
                [0:MAX_VALUE_32 - 1] :/ 2, 
                MAX_VALUE_32 - 1 :/ 2};
    }

    //------------------------------------------------------------------------------
    // The constructor for the sequence.
    //------------------------------------------------------------------------------
    function new(string name ="pc_seq");
        super.new(name);
    endfunction : new

    //------------------------------------------------------------------------------
    // The main task to be executed within the sequence.
    //------------------------------------------------------------------------------
    task body();
        // Create sequence
        req = pc_seq_item::type_id::create("req");
        // Wait for sequencer ready
        start_item(req);
        // Randomize sequence item
        if (!(req.randomize() with {
            req.pc == local::pc;
        })) `uvm_fatal(get_name(), "Failed to randomize")
        // Send to sequencer
        finish_item(req);
        // Wait until request is completed
        get_response(rsp, req.get_transaction_id());
    endtask : body

endclass : pc_seq