//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
interface data2_if ();
    // data2 output signal.
    logic[31:0] data2;
endinterface : data2_if

