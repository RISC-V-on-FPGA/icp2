//------------------------------------------------------------------------------
// control_in_if interface
//
// This interface provides a control_in output signal.
// 
//------------------------------------------------------------------------------
interface control_in_if ();
    // control_in output signal.                    kanske behöver importera komponenter från kommon för att han skall fatta vad control_type är?????????????????????
    control_type control_in;
endinterface : control_in_if

