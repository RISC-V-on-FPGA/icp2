//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
interface ex_mem_RegWrite_if (input logic clk, input logic rst_n);
    // ex_mem_RegWrite output signal.
    logic[31:0] ex_mem_RegWrite;
endinterface : ex_mem_RegWrite_if

