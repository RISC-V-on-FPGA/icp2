//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
interface data1_if (input logic clk, input logic rst_n);
    // data1 output signal.
    logic[31:0] data1;
endinterface : data1_if

