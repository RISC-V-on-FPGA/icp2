//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
interface data1_if ();
    // data1 output signal.
    logic[31:0] data1;
endinterface : data1_if

