//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
interface immediate_data_if ();
    // immediate_data output signal.
    logic[31:0] immediate_data;
endinterface : immediate_data_if

