//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
interface data2_if (input logic clk, input logic rst_n);
    // data2 output signal.
    logic[31:0] data2;
endinterface : data2_if

